module decode (logic input [13:0] opcode);

endmodule //decode
