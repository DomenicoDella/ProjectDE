module decode ();

endmodule //decode
